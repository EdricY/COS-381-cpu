LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE work.p.all;

ENTITY test_b_shifter IS
END test_b_shifter;


ARCHITECTURE test OF test_b_shifter IS
    SIGNAL a, res: word;
    SIGNAL shift_amt: reg_address;
    SIGNAL right_shift, zfl, cfl, ofl, nfl: STD_LOGIC;
BEGIN
    b_shift: ENTITY work.b_shifter(logic) PORT MAP (a, shift_amt, right_shift, res, zfl, cfl, ofl, nfl);


    PROCESS
        TYPE pattern_type IS RECORD
            a: word;
            shift_amt: reg_address;
            right_shift: STD_LOGIC;
            res: word;
            zfl, cfl, ofl, nfl: STD_LOGIC;
        END RECORD;

        TYPE pattern_array IS ARRAY (NATURAL RANGE <>) OF pattern_type;

        CONSTANT patterns: pattern_array :=
            --  a            shift    r     res         z    c    o    n
            ( (x"00000000", "00000", '0', x"00000000", '1', '0', '0', '0'),
              (x"00000007", "00001", '0', x"0000000E", '0', '0', '0', '0'),
              (x"00000007", "00010", '0', x"0000001C", '0', '0', '0', '0'),
              (x"00000007", "00000", '0', x"00000007", '0', '0', '0', '0'),
              (x"00000007", "00100", '0', x"00000070", '0', '0', '0', '0'),
              (x"00000007", "01000", '0', x"00000700", '0', '0', '0', '0'),
              (x"00000007", "10000", '0', x"00070000", '0', '0', '0', '0'),
              (x"00000007", "10100", '0', x"00700000", '0', '0', '0', '0'), 
              (x"00000007", "11000", '0', x"07000000", '0', '0', '0', '0'),
              (x"00000007", "11100", '0', x"70000000", '0', '0', '0', '0'),
              (x"00000007", "11101", '0', x"E0000000", '0', '0', '0', '1'),
              (x"00000007", "11110", '0', x"C0000000", '0', '1', '1', '1'),
              (x"00000007", "11111", '0', x"80000000", '0', '1', '1', '1'),
              (x"FFFFFFFF", "11111", '0', x"80000000", '0', '1', '1', '1'),
              (x"FFFFFFFD", "11111", '0', x"80000000", '0', '0', '1', '1'),
              (x"FFFFFFFC", "11111", '0', x"00000000", '1', '0', '1', '0'), --16

              (x"12345678", "00100", '0', x"23456780", '0', '1', '1', '0'),
              (x"12345678", "10000", '0', x"56780000", '0', '0', '1', '0'),
              (x"12345678", "00100", '1', x"01234567", '0', '1', '1', '0'),
              (x"12345678", "10000", '1', x"00001234", '0', '0', '1', '0'),

              (x"80000000", "10000", '0', x"00000000", '1', '0', '1', '0'),
              (x"80000000", "11111", '1', x"00000001", '0', '0', '0', '0'),
              (x"00008000", "10000", '0', x"80000000", '0', '0', '0', '1'),

              (x"00010000", "10000", '0', x"00000000", '1', '1', '1', '0'),
              (x"01000000", "01000", '0', x"00000000", '1', '1', '1', '0'),
              (x"10000000", "00100", '0', x"00000000", '1', '1', '1', '0'),
              (x"40000000", "00010", '0', x"00000000", '1', '1', '1', '0'),
              (x"80000000", "00001", '0', x"00000000", '1', '1', '1', '0'),

              (x"00018000", "10000", '0', x"80000000", '0', '1', '1', '1'),
              (x"01800000", "01000", '0', x"80000000", '0', '1', '1', '1'),
              (x"18000000", "00100", '0', x"80000000", '0', '1', '1', '1'),
              (x"60000000", "00010", '0', x"80000000", '0', '1', '1', '1'),
              (x"C0000000", "00001", '0', x"80000000", '0', '1', '1', '1'),

              (x"00000000", "00000", '1', x"00000000", '1', '0', '0', '0'),
              (x"E0000000", "00001", '1', x"70000000", '0', '0', '0', '0'),
              (x"E0000000", "00010", '1', x"38000000", '0', '0', '0', '0'),
              (x"E0000000", "00000", '1', x"E0000000", '0', '0', '0', '1'),
              (x"E0000000", "00100", '1', x"0E000000", '0', '0', '0', '0'),
              (x"E0000000", "01000", '1', x"00E00000", '0', '0', '0', '0'),
              (x"E0000000", "10000", '1', x"0000E000", '0', '0', '0', '0'),
              (x"E0000000", "10100", '1', x"00000E00", '0', '0', '0', '0'),
              (x"E0000000", "11000", '1', x"000000E0", '0', '0', '0', '0'),
              (x"E0000000", "11100", '1', x"0000000E", '0', '0', '0', '0'),
              (x"E0000000", "11101", '1', x"00000007", '0', '0', '0', '0'),
              (x"E0000000", "11110", '1', x"00000003", '0', '1', '1', '0'),
              (x"E0000000", "11111", '1', x"00000001", '0', '1', '1', '0'),
              (x"FFFFFFFF", "11111", '1', x"00000001", '0', '1', '1', '0'),
              (x"BFFFFFFF", "11111", '1', x"00000001", '0', '0', '1', '0'),
              (x"3FFFFFFF", "11111", '1', x"00000000", '1', '0', '1', '0'),

              (x"00000000", "00000", '1', x"00000000", '1', '0', '0', '0')
            );
    
    BEGIN
        FOR i IN patterns'range LOOP
            a <= patterns(i).a;
            shift_amt <= patterns(i).shift_amt;
            right_shift <= patterns(i).right_shift;

            wait for 1 ms;

            assert res = patterns(i).res
                report "bad result" severity error;
            assert zfl = patterns(i).zfl
                report "bad zfl" severity error;
            assert cfl = patterns(i).cfl
                report "bad cfl" severity error;
            assert ofl = patterns(i).ofl
                report "bad ofl" severity error;
            assert nfl = patterns(i).nfl
                report "bad nfl" severity error;
        END LOOP;

        assert false
            report "end of b_shifter test" severity note;

        wait;
    END PROCESS;
END test;
